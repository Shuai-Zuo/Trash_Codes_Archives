module functout(state,opcode,funct,zero,PCWr,IRWr,MemtoReg,RegWr,ALUsrc,MemWr,Extop,RegDst,npc_sel,ALUctr,sbsel,lbsel);
input [3:0]state;
input [5:0]opcode,funct;
input zero;
output reg PCWr,IRWr,ALUsrc,MemWr,RegWr,Extop,sbsel,lbsel;
output reg [2:0]npc_sel;
output reg [1:0]MemtoReg,RegDst;
output reg [2:0]ALUctr;
parameter [3:0]IF = 4'b0000, 
               ID = 4'b0001,
               MA = 4'b0010,
               MR = 4'b0011,
               MemWB = 4'b0100,
               MW = 4'b0101,
               Exe = 4'b0110,
               WB = 4'b0111,
               Branch = 4'b1000,
               Jump = 4'b1001;
               parameter [5:0]R=6'b000000,
                              addu=6'b100001,
                              subu=6'b100011,
                              slt=6'b101010,
                              jr=6'b001000,
                              addi=6'b001000,
                              addiu=6'b001001,
                              ori=6'b001101,
                              lui=6'b001111,
                              sw=6'b101011,
                              lw=6'b100011,
                              sb=6'b101000,
                              lb=6'b100000,
                              beq=6'b000100,
                              j=6'b000010,
                              jal=6'b000011,
                              jalr=6'b001001;
 always@(state)
 begin
   if(state==IF||state==Jump) PCWr=1;
   else PCWr=0;
     
   if(state==IF) IRWr=1;
   else IRWr=0;
     
   if(state==MA) 
     if(opcode==sw||opcode==sb) MemWr=1;
     else MemWr=0;
   else MemWr=0;
     
   if(state==MemWB||state==WB||(opcode==jal && state==Jump)||(funct==jalr && state == Jump))
     RegWr=1;
   else RegWr=0;
     
   case(opcode)
     R:begin
       case(funct)
         addu:begin npc_sel=3'b000;RegDst=2'b01;ALUsrc=0;MemtoReg=2'b00;ALUctr=3'b000;end
         subu:begin npc_sel=3'b000;RegDst=2'b01;ALUsrc=0;MemtoReg=2'b00;ALUctr=3'b001;end
         slt:begin npc_sel=3'b000;RegDst=2'b01;ALUsrc=0;MemtoReg=2'b00;ALUctr=3'b100;end
         jr:begin npc_sel=3'b011;end
       endcase
       end
         addi :begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b00;ALUctr=3'b000;Extop=1;end
         addiu:begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b00;ALUctr=3'b000;Extop=1;end
         ori:  begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b00;ALUctr=3'b010;Extop=0;end
         lui:  begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b00;ALUctr=3'b011;Extop=0;end
         sw:   begin npc_sel=3'b000;ALUsrc=1;ALUctr=3'b000;Extop=1;sbsel=0;end
         lw:   begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b01;ALUctr=3'b000;Extop=1;lbsel=0;end
         sb:   begin npc_sel=3'b000;ALUsrc=1;ALUctr=3'b000;Extop=1;sbsel=1;end
         lb:   begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=1;MemtoReg=2'b01;ALUctr=3'b000;Extop=1;lbsel=1;end
         beq:  begin 
               ALUctr=3'b001;
               if(zero)npc_sel=3'b001;
               else npc_sel=3'b000;
               end
         j:npc_sel=3'b010;
         jal:begin npc_sel=3'b010;RegDst=2'b10;MemtoReg=2'b10;end
         
         default: begin npc_sel=3'b000;RegDst=2'b00;ALUsrc=0;MemtoReg=2'b00;ALUctr=3'b000;Extop=0;sbsel=0;lbsel=0;end
    endcase
 end
endmodule