library verilog;
use verilog.vl_types.all;
entity exp9_vlg_vec_tst is
end exp9_vlg_vec_tst;
