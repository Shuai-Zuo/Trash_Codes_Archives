library verilog;
use verilog.vl_types.all;
entity data_deal_vlg_vec_tst is
end data_deal_vlg_vec_tst;
