library verilog;
use verilog.vl_types.all;
entity nambscld_vlg_vec_tst is
end nambscld_vlg_vec_tst;
