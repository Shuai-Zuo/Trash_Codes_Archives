module scan2(CLK,SEL,QA,QB,QC,QD,QE,QF,QG,QH);
input CLK;
output[2:0]SEL;
reg[2:0]SEL;
output QA,QB,QC,QD,QE,QF,QG,QH;
reg QA,QB,QC,QD,QE,QF,QG,QH;
always@(posedge CLK)
begin
	case(SEL)
		3'b000:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11111101;
		3'b001:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11111011;
		3'b010:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11110111;
		3'b011:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11101111;
		3'b100:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11011111;
		3'b101:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b10111111;
		3'b110:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b01111111;
		3'b111:{QH,QG,QF,QE,QD,QC,QB,QA}<=8'b11111110;
	endcase
	SEL<=SEL+1'b1;
end
endmodule