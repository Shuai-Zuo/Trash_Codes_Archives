library verilog;
use verilog.vl_types.all;
entity exp_5_vlg_tst is
end exp_5_vlg_tst;
