library verilog;
use verilog.vl_types.all;
entity IR is
    port(
        clk             : in     vl_logic;
        IRWr            : in     vl_logic;
        IR_in           : in     vl_logic_vector(31 downto 0);
        opcode          : out    vl_logic_vector(5 downto 0);
        rs              : out    vl_logic_vector(4 downto 0);
        rt              : out    vl_logic_vector(4 downto 0);
        rd              : out    vl_logic_vector(4 downto 0);
        imm             : out    vl_logic_vector(15 downto 0);
        funct           : out    vl_logic_vector(5 downto 0);
        \IMM\           : out    vl_logic_vector(25 downto 0)
    );
end IR;
