library verilog;
use verilog.vl_types.all;
entity selection_vlg_vec_tst is
end selection_vlg_vec_tst;
