library verilog;
use verilog.vl_types.all;
entity redw_vlg_vec_tst is
end redw_vlg_vec_tst;
