library verilog;
use verilog.vl_types.all;
entity controlltst_vlg_vec_tst is
end controlltst_vlg_vec_tst;
