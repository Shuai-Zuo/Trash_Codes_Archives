module dm_1k(addr,din,dout,we,sbsel);
  input [31:0] din;
  input [9:0] addr;
  input we,sbsel;
  output [31:0] dout;
  //reg [31:0] dout;
  reg [7:0] dm[1023:0];
  integer i;
  //assign sw_addr=addr[9:0];
  //assign sb_addr=addr[1:0];
  initial
  begin
    for(i=0;i<1024;i=i+1)
      dm[i]=0;
  end
  always@(we) //addr or or din or sbsel 
  begin
    if(we==1'b1)
      begin
        if(sbsel)
          begin
            dm[addr]=din[7:0];
          end
        else   
        begin
          dm[addr]=din[7:0];
          dm[addr+1]=din[15:8];
          dm[addr+2]=din[23:16];
          dm[addr+3]=din[31:24];
        end
      end
    
  end
    //always@(addr or we or din)
    //begin
     // if(we==1'b0)
     //   dout={dm[addr[9:0]+3],dm[addr[9:0]+2],dm[addr[9:0]+1],dm[addr[9:0]]};
    //end
    assign dout={dm[addr+3],dm[addr+2],dm[addr+1],dm[addr]};
endmodule
  
