library verilog;
use verilog.vl_types.all;
entity exp6_top_vlg_vec_tst is
end exp6_top_vlg_vec_tst;
