library verilog;
use verilog.vl_types.all;
entity controlltst_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        result_Con      : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end controlltst_vlg_sample_tst;
