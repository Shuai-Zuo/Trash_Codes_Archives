library verilog;
use verilog.vl_types.all;
entity a31_vlg_vec_tst is
end a31_vlg_vec_tst;
