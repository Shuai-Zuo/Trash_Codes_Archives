library verilog;
use verilog.vl_types.all;
entity e11_vlg_vec_tst is
end e11_vlg_vec_tst;
