module control(clk,reset,result_Con,consignal,sel_Con,inc_Floor,red_Floor,ce,up_d,stop_r,rst,ce_Count,state);
parameter S0=4'b0000,S1=4'b0001,S2=4'b0010,S3=4'b0011,S4=4'b0100,S5=4'b0101,S6=4'b0110,S7=4'b0111,S8=4'b1000,S9=4'b1001,S10=4'b1010,S11=4'b1011,S12=4'b1100,S13=4'b1101,S14=4'b1110,S15=4'b1111;
input clk,reset,result_Con,consignal;
  output [1:0] sel_Con;
  output inc_Floor,red_Floor,ce,up_d,stop_r,rst,ce_Count;
  output [3:0]state;
  reg [1:0] sel_Con;
  reg inc_Floor,red_Floor,ce,up_d,stop_r,rst,ce_Count;
  reg[3:0] state;
always @ (posedge clk or negedge reset)
  begin
   if(!reset)
   state<=S0;
  else
  begin
   case(state)
   S0:state<=S1;
   S1:if(result_Con)
    state<=S3;
    else
    state<=S2;
   S2:if(result_Con)
    state<=S9;
    else
    state<=S1;
   S3:state<=S4;
   S4:if(consignal)
    begin
    state<=S5;
    end
      else
   state<=S4;
   S5:state<=S6;
   S6:if(result_Con)
	state<=S8;
	else
	state<=S7;
   S7:if(result_Con)
	state<=S4;
	else
	state<=S8;
   S8:if(consignal)
	begin
	state<=S1;
	end
	else
	state<=S8;
   S9:state<=S10;
   S10:if(consignal)
	begin
	state<=S11;
	end
	else
	state<=S10;
   S11:state<=S12;
   S12:if(result_Con)
	state<=S14;
	else
	state<=S13;
   S13:if(result_Con)
	state<=S10;
	else
	state<=S14;
   S14:if(consignal)
	begin
	state<=S2;
	end
	else
	state<=S14;
   default:state<=S15;
   endcase
   end
end
	always @ (state)  
	begin
	case(state)
	S0:
	begin
	rst=1;
	red_Floor<=0;
	inc_Floor<=0;
	stop_r<=0;
	up_d<=0;
	ce<=0;
	end
	S1: 
	begin
   ce<=1;
   rst<=0;
   ce_Count<=0;
   sel_Con<=2'b00;
   end
	S2:
	begin
   ce<=1;
	rst<=0;
   ce_Count<=0;
   sel_Con<=2'b01;
   end
	S3:
	begin
   up_d<=0;
	rst<=0;
   stop_r<=1;
   ce<=0;
   end
	S4:
	begin
   ce_Count<=1;
	rst<=0;
   end
	S5:
	begin
   ce_Count<=0;
	rst<=0;
   inc_Floor<=1;
   end
	S6:
	begin
   inc_Floor<=0;
	rst<=0;
   sel_Con<=2'b10;
   end
	S7:
	begin
   sel_Con<=2'b00;
	rst<=0;
   end
	S8:
	begin
   ce<=1;
   stop_r<=0;
	rst<=0;
   ce_Count<=1;
   end
	S9:
	begin 
   up_d<=1;
	rst<=0;
   stop_r<=1;
   ce<=0;
   end
	S10:
	begin
	rst<=0;
   ce_Count<=1;
   end
	S11:
	begin
	rst<=0;
   ce_Count<=0;
	red_Floor<=1;
   end
   S12:
	begin
	rst<=0;
   red_Floor<=0;
   sel_Con<=2'b11;
   end
	S13:
	begin
	rst<=0;
   sel_Con<=2'b01;
	end
	S14:
	begin
	rst<=0;
   ce<=1;
   stop_r<=0;
   ce_Count<=1;
   end
	//default:state<=S15;
	endcase
   end
endmodule

