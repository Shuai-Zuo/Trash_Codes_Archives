library verilog;
use verilog.vl_types.all;
entity exp6_vlg_tst is
end exp6_vlg_tst;
