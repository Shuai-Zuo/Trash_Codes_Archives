library verilog;
use verilog.vl_types.all;
entity experiment31_vlg_vec_tst is
end experiment31_vlg_vec_tst;
