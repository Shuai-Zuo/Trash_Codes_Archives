module Extender(ExtOp,imm,imm_out);
  input ExtOp;
  input[15:0] imm;
  output [31:0] imm_out;
  reg[31:0] imm_out;
  
  always@(imm or ExtOp)
  begin
    if(!ExtOp)
      imm_out = {{16{1'b0}},imm[15:0]};
    else
      imm_out = {{16{imm[15]}},imm[15:0]};
  end
endmodule
