library verilog;
use verilog.vl_types.all;
entity exp8_top_vlg_vec_tst is
end exp8_top_vlg_vec_tst;
