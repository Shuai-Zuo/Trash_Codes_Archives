library verilog;
use verilog.vl_types.all;
entity condition_vlg_vec_tst is
end condition_vlg_vec_tst;
