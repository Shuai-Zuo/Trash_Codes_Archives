library verilog;
use verilog.vl_types.all;
entity t2_vlg_vec_tst is
end t2_vlg_vec_tst;
