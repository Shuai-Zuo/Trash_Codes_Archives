library verilog;
use verilog.vl_types.all;
entity exp10_vlg_vec_tst is
end exp10_vlg_vec_tst;
