/*module move(in1,in2,in3,in4,in5,in6,in7,in8,pressed,key,out1,out2,out3,out4,out5,out6,out7,out8);
input[3:0]in1,in2,in3,in4,in5,in6,in7,in8;
input pressed;
input[3:0]key;
output[3:0]out1,out2,out3,out4,out5,out6,out7,out8;
always@(posedge pressed)
begin
{out1,out2,out3,out4,out5,out6,out7,out8}<={key,in1,in2,in3,in4,in5,in6,in7};
end
endmodule*/