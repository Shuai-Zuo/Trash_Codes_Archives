library verilog;
use verilog.vl_types.all;
entity indoor_request_vlg_vec_tst is
end indoor_request_vlg_vec_tst;
