library verilog;
use verilog.vl_types.all;
entity red_vlg_vec_tst is
end red_vlg_vec_tst;
