library verilog;
use verilog.vl_types.all;
entity keyboard_scan_vlg_vec_tst is
end keyboard_scan_vlg_vec_tst;
