library verilog;
use verilog.vl_types.all;
entity counter_vlg_check_tst is
    port(
        con             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end counter_vlg_check_tst;
