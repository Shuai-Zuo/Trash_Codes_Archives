library verilog;
use verilog.vl_types.all;
entity scan_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end scan_vlg_sample_tst;
