library verilog;
use verilog.vl_types.all;
entity experimentIII_vlg_vec_tst is
end experimentIII_vlg_vec_tst;
