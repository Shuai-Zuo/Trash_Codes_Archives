module condition(get_dest,get_call,cur_Floor,sel_condition,clk,result);
input [3:0]get_dest;
input [5:0]get_call;
input [1:0]sel_condition;
input clk;
input [1:0]cur_Floor;
output result;
reg result;
integer flag,i;
always@(posedge clk)
begin
case(sel_condition)
2'b00:
begin
case(cur_Floor)
2'b00:
begin
if(get_dest[1]||get_dest[2]||get_dest[3]||get_call[1]||get_call[2]||get_call[3]||get_call[4]||get_call[5])
	result=1;
else
	result=0;
end
2'b01:
begin
if(get_dest[2]||get_dest[3]||get_call[3]||get_call[4]||get_call[5])
	result=1;
else
	result=0;
end
2'b10:
begin
if(get_dest[3]||get_call[5])
	result=1;
else
	result=0;
end
default:result=0;
endcase
end
2'b01:
begin
case(cur_Floor)
2'b11:
begin
if(get_dest[0]||get_dest[1]||get_dest[2]||get_call[0]||get_call[2]||get_call[4])
	result=1;
else
	result=0;
end
2'b10:
begin
if(get_dest[0]||get_dest[1]||get_call[0]||get_call[2])
	result=1;
else
	result=0;
end
2'b01:
begin
if(get_dest[0]||get_call[0])
	result=1;
else
	result=0;
end
default:result=0;
endcase
end
2'b10:
begin
case(cur_Floor)
2'b00:
begin
if(get_dest[0]||get_call[0])
	result=1;
else
	result=0;
end
2'b01:
begin
if(get_dest[1]||get_call[1])
	result=1;
else
	result=0;
end
2'b10:
begin
if(get_dest[2]||get_call[3])
	result=1;
else
	result=0;
end
2'b11:
begin
if(get_dest[3])
	result=1;
else
	result=0;
end
default:result=0;
endcase
end
2'b11:
begin
case(cur_Floor)
2'b00:
begin
if(get_dest[0])
	result=1;
else
	result=0;
end
2'b01:
begin
if(get_dest[1]||get_call[2])
	result=1;
else
	result=0;
end
2'b10:
begin
if(get_dest[2]||get_call[4])
	result=1;
else
	result=0;
end
2'b11:
begin
if(get_dest[3]||get_call[5])
	result=1;
else
	result=0;
end
default:result=0;
endcase
end
endcase
end
endmodule
