module gpr(ReadReg1,ReadReg2,WriteReg,WriteData,ReadData1,ReadData2,RegWrite,rst,OF);
input [4:0] ReadReg1,ReadReg2,WriteReg;
input [31:0] WriteData;
input RegWrite,rst,OF;
output [31:0] ReadData1,ReadData2;
reg [31:0] register[31:0];
integer i;
assign ReadData1=register[ReadReg1];
assign ReadData2=register[ReadReg2];
always @( RegWrite or rst)
begin
  if(rst==1'b1)
    begin
      for(i=0;i<31;i=i+1)
        register[i]=0;
    end
  else
    begin
      if(RegWrite==1'b1 && WriteReg !=5'b00000)
        register[WriteReg]=WriteData;
    end
end
always@(negedge OF)
begin
  register[30]=1;
  register[22]=0;
end
endmodule
