library verilog;
use verilog.vl_types.all;
entity selection_8t1_vlg_vec_tst is
end selection_8t1_vlg_vec_tst;
